module top:
	
endmodule 